----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/22/2021 09:22:50 PM
-- Design Name: 
-- Module Name: controller - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity controller is
--  Port ( );
generic(CCW : INTEGER := 32;
        CCWdiv8 : INTEGER := 4);
port(
     clk, rst: in STD_LOGIC;
    -- INPUT FROM CYRPTO CORE
     bdi_type: in STD_LOGIC_VECTOR(3 downto 0);
     msg_auth_ready, decrypt_in, bdi_eoi, bdi_eot, bdo_ready, key_update, key_valid, bdi_valid: in STD_LOGIC;
     -- SIGNALS GENERATED BY CONTROLLER FOR DATAPATH
     selInitial, selS, selSR, selD, selT: out STD_LOGIC;
     enRound, enTK, enKey, enAM, enN, enS, enDD, enCI_T: out STD_LOGIC;
     Bin : STD_LOGIC_VECTOR(3 downto 0);
     -- OUTPUT for CRYPTO CORE
     end_of_block, bdo_valid, msg_auth, msg_auth_valid, bdi_ready: out STD_LOGIC;
     bdo_type: out STD_LOGIC_VECTOR(3 downto 0);
     bdo_valid_bytes: out STD_LOGIC_VECTOR(CCWdiv8-1 downto 0));
end controller;

architecture Behavioral of controller is

begin


end Behavioral;
