----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/22/2021 09:22:50 PM
-- Design Name: 
-- Module Name: controller - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity controller is
--  Port ( );
generic(CCW : INTEGER := 32;
        CCWdiv8 : INTEGER := 4);
port(
     clk, rst: in STD_LOGIC;
    -- INPUT FROM CYRPTO CORE
     bdi_type: in STD_LOGIC_VECTOR(3 downto 0);
     msg_auth_ready, decrypt_in, bdi_eoi, bdi_eot, bdo_ready, key_update, key_valid, bdi_valid: in STD_LOGIC;
     -- INPUT FROM DATAPATH
     tag_verify : in STD_LOGIC;
     E_done : in STD_LOGIC;
     -- SIGNALS GENERATED BY CONTROLLER FOR DATAPATH
     E_start : out STD_LOGIC;
     selS, selSR, selD, selT, selMR: out STD_LOGIC;
     selAM : out STD_LOGIC_VECTOR(1 downto 0);
     enKey, enAM, enN, enS, enDD, enCI_T, enTag: out STD_LOGIC;
     Bin :out STD_LOGIC_VECTOR(4 downto 0);
     ldCi_T : out STD_LOGIC;
     Len8 : out STD_LOGIC_VECTOR(7 downto 0);
     -- OUTPUT for CRYPTO CORE
     end_of_block, bdo_valid, msg_auth, msg_auth_valid, bdi_ready, key_ready: out STD_LOGIC;
     bdo_type: out STD_LOGIC_VECTOR(3 downto 0);
     bdo_valid_bytes: out STD_LOGIC_VECTOR(CCWdiv8-1 downto 0));
end controller;

architecture Behavioral of controller is
type state is (idle, load_key, load_npub, wait_ad, load_ad, pad_ad, rho_ad, ek_ad, rho_ad_pad, ek_ad_pad, rho_final, ek_nonce, load_data, process_tag, output_tag, verify_tag);
signal state_reg, state_next : state;

-- register to store bdi_valid bytes and output for when output of Data is passed through
signal bdi_vb_reg : std_logic_vector(15 downto 0);
signal bdi_vb_reg_next : std_logic_vector(3 downto 0);
signal envb : std_logic;

signal numB_s_next, numB_s : unsigned(55 downto 0);
signal numB_s_vec : std_logic_vector(55 downto 0);

signal len8_s_next, len8_s : unsigned(7 downto 0);

signal cnt_s_next, cnt_s : integer range 0 to 4;

-- Constants for bdi/bdo type encodings

constant HDR_AD : std_logic_vector(3 downto 0) := "0001";
constant HDR_PT : std_logic_vector(3 downto 0) := "0100";
constant HDR_CT : std_logic_vector(3 downto 0) := "0101";
constant HDR_TAG : std_logic_vector(3 downto 0) := "1000";
constant HDR_KEY : std_logic_vector(3 downto 0) := "1100";
constant HDR_NPUB : std_logic_vector(3 downto 0) := "1101";
constant HDR_HASH_MSG : std_logic_vector(3 downto 0) := "0111";
constant HDR_HASH_VALUE : std_logic_vector(3 downto 0) := "1001";

-- internal flags
signal pad_block_status : std_logic;

begin
-- raw connections
numB_s_vec <= std_logic_vector(numB_s);

Len8 <= std_logic_vector(len8_s);


-- process reg for storing bdi_type for message
process(clk)
begin
    if rising_edge(clk) then
        if envb = '1' then
            bdi_vb_reg <= bdi_vb_reg(11 downto 0) & bdi_vb_reg_next;
        end if;
    end if;    
end process;


-- state register
process(clk)
begin
    if rising_edge(clk) then
        if rst = '1' then
            state_reg <= idle;
            pad_block_status <= '0';
            cnt_s <= 0;
            numB_s <= (others => '0');
            cnt_s <= 0;
            pad_block_status <= '0';
        else
            state_reg <= state_next;
            cnt_s <= cnt_s_next;
            numB_s <= numB_s_next;
            
        end if;
    end if;
end process;


-- next state register
process(state_reg, key_valid, bdi_valid, bdi_eoi, bdo_ready, bdi_eot, cnt_s, bdi_vb_reg, decrypt_in, len8_s, E_done, numB_s_vec, numB_s, bdi_type)
    begin
    
    cnt_s_next <= cnt_s;
    bdi_vb_reg_next <= (others => '0');
    key_ready <= '0';
    Bin <= (others => '0');
    enDD <= '0';
    selS <= '0';
    selSR <= '0';
    enS <= '0';
    selT <= '0';
    selD <= '0';
    enKey <= '0';
    
    case state_reg is
        
        when idle =>
            if key_valid = '1' then
                if key_update = '1' then
                    state_next <= load_key;
                elsif bdi_valid = '1' then
                    state_next <= load_npub;
                else 
                    state_next <= idle;
                end if;
            elsif bdi_valid = '1' then
                state_next <= load_npub;
            else 
                state_next <= idle;
            end if;
         
         when load_key =>
                key_ready <= '1';        
                if key_valid = '0' then
                    state_next <= load_key;
                elsif cnt_s = 4 then
                    cnt_s_next <= 0;
                    state_next <= idle;
                else 
                    cnt_s_next <= cnt_s + 1;
                    enKey <= '1';
                    state_next <= load_key;
                end if;
                
         when load_npub =>
                bdi_ready <= '1';
                if bdi_valid = '1' then
                    if bdi_type = HDR_NPUB then
                        if cnt_s = 4 then
                            cnt_s_next <= 0;
                            if bdi_eoi = '1' then
                                state_next <= process_tag;
                                -- need to look at this segment of code more closely
                            else 
                                state_next <= wait_ad;
                            end if;
                        else
                            cnt_s_next <= cnt_s + 1;
                            enN <= '1';
                            state_next <= load_npub;
                        end if;
                    else
                        state_next <= load_npub;
                    end if;
                else
                    state_next <= load_npub;
                end if;
                
         when wait_ad =>
                if bdi_type = HDR_AD then
                    numB_s_next <= (others => '0');
                    state_next <= load_ad;
                else
                    state_next <= load_data;
                end if;
                    
         when load_ad =>
                bdi_ready <= '1';
                if bdi_valid = '0' then
                    state_next <= load_ad;
                else
                    if cnt_s = 4 then
                        pad_block_status <= '0';
                        cnt_s_next <= 0;
                        numB_s_next <= numB_s + 1;
                        if numB_s_vec(0) = '1' then
                            state_next <= ek_ad;
                        else 
                            state_next <= rho_ad;
                        end if;
                    else
                        if bdi_eot = '1' then 
                            cnt_s_next <= cnt_s + 1;
                            enAM <= '1';
                            pad_block_status <= '1';
                            state_next <= pad_ad;
                        else
                            cnt_s_next <= cnt_s + 1;
                            enAM <= '1';
                            state_next <= load_ad;
                        end if;
                    end if;
                end if;
             
              -- Did not get to implement the rest of the main controller in vhdl
              
         when pad_ad =>
                if cnt_s < 3 then
                    cnt_s_next <= cnt_s + 1;
                    selAM <= "01";
                    state_next <= pad_ad;
                else
                    if cnt_s = 4 then
                        cnt_s_next <= 0;
                        numB_s_next <= numB_s + 1;
                        if numB_S(0) = '1' then
                            state_next <= ek_ad_pad;
                        else
                            state_next <= rho_ad_pad;
                        end if;
                    else
                        cnt_s_next <= cnt_s + 1;
                        selAM <= "10";
                        state_next <= pad_ad;
                    end if;
                end if;
            
         when ek_ad =>
                E_start <= '1';
                Bin <= "01000";                                            
                if E_done = '1' then
                    enDD <= '1';
                    state_next <= load_ad;
                else
                    selS <= '1';
                    state_next <= ek_ad;
                end if;
         
         when rho_ad =>
                if numB_S_vec = x"00000000000001" then
                    selSR <= '1';
                    enS <= '1';
                    state_next <= load_ad;
                else
                    enDD <= '1';
                    enS <= '1';
                    state_next <= load_ad;
                end if;
         
         when rho_ad_pad =>
                if numB_S_vec = x"00000000000001" then
                    selSR <= '1';
                    enS <= '1';
                    enDD <= '1';
                    state_next <= rho_final;
                else
                    enS <= '1';
                    enDD <= '1';
                end if;
         
         when ek_ad_pad =>
                E_start <= '1';
                Bin <= "01000";                                            
                if E_done = '1' then
                    selMR <= '1';
                    enS <= '1';
                    state_next <= rho_final;
                else 
                    state_next <= ek_ad_pad;
                end if;
         
         when rho_final =>
                if len8_s = x"FF" then
                    E_start <= '1';
                    Bin <= "11000";
                    selT <= '1';
                    state_next <= ek_nonce;
                else
                    E_start <= '1';
                    Bin <= "11010";
                    selT <= '1';
                    state_next <= ek_nonce;
                end if;
         
         when ek_nonce =>
                 if E_done = '1' then
                    selD <= '1';
                    enDD <= '1';
                    state_next <= load_data;
                 else
                    state_next <= ek_nonce;
                 end if;
         
         when load_data =>
                bdi_ready <= '1';
                if bdi_valid = '1' then
                    if cnt_s = 4 then
                        pad_block_status <= '1';
                        cnt_s_next <= 0;
                        numB_s_next <= numB_s + 1;
                    -- else
                       -- if bdi_eot = '1' then
                    end if;
                end if;
                            -- ran out of time to implement but it is very similiar to what should occur during Loading of Message just now cipher input is Nonce
                            -- and some small very miniscule other changes are to be expected.
            -- After this, subsequent changes would be made in order to effectively Process each method into Rho Function or TBC call, and corresponding output would
            -- fed into the PISO for loading data out through bdo port. We also compare data that is stored with loaded tag later on in last TBC and Rho function call in order
            -- to verify that the two tags are exactly the same for message authentication purposes
         
         when process_tag =>
                if cnt_s = 4 then
                    cnt_s_next <= 0;
                    if decrypt_in = '1' then
                        state_next <= verify_tag;
                    else
                        state_next <= output_tag;
                    end if;
                else
                    cnt_s_next <= cnt_s + 1;
                    enTag <= '1';
                end if;
                     
         when verify_tag =>
                bdi_ready <= '1';
                
         when output_tag =>
                cnt_s_next <= cnt_s;
    end case;
    
end process;



end Behavioral;
